module UART_TOP(TX_IN_P, TX_IN_V, PAR_EN, PAR_TYP, TX_CLK, RST, RX_CLK, Prescale, RX_OUT_V, RX_OUT_P, TX_OUT_S, TX_OUT_V);
parameter WIDTH = 8, START_BIT = 0, STOP_BIT = 1;
input [WIDTH-1:0] TX_IN_P;
input TX_IN_V, PAR_EN, PAR_TYP, TX_CLK, RST, RX_CLK;
input [8:0] Prescale;
output TX_OUT_S, TX_OUT_V;
output [WIDTH-1:0] RX_OUT_P;
output RX_OUT_V;
UART_TX#(WIDTH,START_BIT,STOP_BIT) TX (TX_IN_P,TX_IN_V,PAR_EN,PAR_TYP,TX_CLK,RST,TX_OUT_S,TX_OUT_V);
UART_RX#(WIDTH,START_BIT,STOP_BIT) RX (TX_OUT_S,Prescale,PAR_EN,PAR_TYP,RST,RX_CLK,RX_OUT_V,RX_OUT_P);
endmodule